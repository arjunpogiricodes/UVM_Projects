







// destination transaction class

class destin_xtn extends uvm_sequence_item;


// factory registration

       `uvm_object_utils(destin_xtn)

// declare the rand feilds



// declare the constructions



// fcuntion new constructor


        function new(string name = "destin_xtn");

                 super.new(name);


        endfunction 



endclass
